-- This is a comment


entity main is
end main;

architecture Behavioral of main is
begin
end Behavioral;
